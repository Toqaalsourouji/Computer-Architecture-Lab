module inverter( input signal , output inverted );
assign inverted= ~signal;
endmodule
