module InstructionMem(input [5:0] addr, output [31:0] data_out);
reg [31:0] mem [0:63];

assign data_out = mem[addr];

initial begin

mem[0] =  32'b00000000011000101000001000110011;
mem[1] =  32'b01000001001101100000001110110011;
mem[2] =  32'b00000101000001100000010001100011;
mem[3] =  32'b00000001101110001000000010110011;
mem[4] =  32'b00000000010000101111111110110011;

end
endmodule
